rem   
rem  PERFORM A DISK TO DISK BACKUP OF FOLDERS ON FILE SERVER
rem
F:
rem
CD F:\DATA
COPY *.* C:\SRVRBKUP\DATA\*.*
rem
CD F:\INCLUDES
COPY *.* C:\SRVRBKUP\INCLUDES\*.*
rem
CD F:\INCLUDES.CNV
COPY *.* C:\SRVRBKUP\INCLUDES.CNV\*.*
rem
CD F:\SOURCE
COPY *.* C:\SRVRBKUP\SOURCE\*.*
rem
CD F:\SOURCE.CNV
COPY *.* C:\SRVRBKUP\SOURCE.CNV\*.*
rem
CD F:\PLC
COPY *.* C:\SRVRBKUP\PLC\*.*
rem
CD F:\SUNBELT
COPY *.* C:\SRVRBKUP\SUNBELT\*.*
rem
CD F:\SUNBELT\CODE
COPY *.* C:\SRVRBKUP\SUNBELT\CODE\*.*
rem
CD F:\SUNBELT\DEMO
COPY *.* C:\SRVRBKUP\SUNBELT\DEMO\*.*
rem
CD F:\UTILS
COPY *.* C:\SRVRBKUP\UTILS\*.*
rem
CD F:\UTILS.CNV
COPY *.* C:\SRVRBKUP\UTILS.CNV\*.*
rem
CD F:\BACKUP
COPY *.* C:\SRVRBKUP\BACKUP\*.*
rem
rem
rem
rem    BE SURE TO CHECK THE COPIES AND SEE IF IT WORKED !
rem
C:
CD C:\WINDOWS
EXIT
